module registers(
input [7:0]
);
endmodule
